module main

fn main() {
	mut age := 20
	println(age)
	age = 21
	println(age)
}
