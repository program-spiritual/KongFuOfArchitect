module main
import os
fn main() {
println(os.args)
}


