module main

fn main() {
	mut a := 0
	mut b := 1
	println('${a}, ${b}') // 0, 1
	a, b = b, a
	println('${a}, ${b}') // 1, 0
}
