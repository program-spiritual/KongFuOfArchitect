module error

fn main() {
  a := 10
  if true {
    a := 20 // error: redefinition of `a`
  }
  // warning: unused variable `a`
}
