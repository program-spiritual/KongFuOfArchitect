module main

a := 0x7B
b := 0b01111011
c := 0o173
println(a)
println(b)
println(c)
num := 1_000_000 // same as 1000000
three := 0b0_11 // same as 0b11
float_num := 3_122.55 // same as 3122.55
hexa := 0xF_F // same as 255
oct := 0o17_3 // same as 0o173
println(num)
println(three)
println(float_num)
println(hexa)
println(oct)
println('/n next line :')
a1 := i64(123)
b1 := u8(42)
c1 := i16(12345)
println(a1)
println(b1)
println(c1)
