module main

for i := 0; i < 10; i++ {
	if i == 6 {
		continue
	}
	print(i)
}
