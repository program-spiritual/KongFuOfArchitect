module main

my_int := 1

my_closure := fn [my_int] () {
	println(my_int)
}

my_closure()
